`timescale 1ns / 1ps

module SN54LS153 (
// port list
	o_1Y	, // output 
	o_2Y	, 
	i_B		, // select
	i_A		, 
	i_1G	, // strobe(active low)
	i_2G	, 
	i_1C0	, // input for o_1Y
	i_1C1	, 
	i_1C2	, 
	i_1C3	, 
	i_2C0	, // input for o_2Y 
	i_2C1	, 
	i_2C2	, 
	i_2C3


);
// port declaration
output 	o_1Y		;
output 	o_2Y		;
input 	i_B			;
input 	i_A			;
input 	i_1G		;
input 	i_2G		;
input 	i_1C0		;
input 	i_1C1		;
input 	i_1C2		;
input 	i_1C3		;
input 	i_2C0		;
input 	i_2C1		;
input 	i_2C2		;
input 	i_2C3		;


// EXAM: behavioral modeling 




endmodule
